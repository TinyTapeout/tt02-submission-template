// Tiny Tapeout 02
// Verilog Template
//Note: available cells can be found in /src/cells.v
//you can also implicitly declare cells using verilog syntax:
//e.g. reg example_dff;
//e.g. assign io_out[2] = usersignal & !dff_q;

module githubusername_top_template(	  //prepend your github username to the top module
	input  [7:0] io_in,		              //do not change port names 
	output [7:0] io_out);
	

 	//*********** Your Design Below ************


endmodule
