// TinyTapeout02: Verilog Template
// Remember to include your top module name in the info.yaml file

module githubusername_top( //prepend your github username
	input  [7:0] io_in,    //leave the port names unchanged
	output [7:0] io_out);

	//****Your Design Here****

endmodule
