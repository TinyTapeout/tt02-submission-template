module toplevel();
endmodule
