// TinyTapeout02: Verilog Template
// Remember to include your top module name in the info.yaml file
// Note: available cells can be found in /src/cells.v
// you can also implicitly declare cells using verilog syntax:
// e.g. reg example_dff;
// e.g. assign io_out[2] = usersignal & !dff_q;

module githubusername_top( //prepend your github username
	input  [7:0] io_in,    //leave the port names unchanged
	output [7:0] io_out);

	//****Your Design Here****

endmodule
